[aimspice]
[description]
213
INVERSOR SIMPLU ANALIZA SEMNAL PULSE
R1 in 1 1k
Rc out ec 1k
C1 in 1 30p
Q out 1 0 Tranzistor
C2 out 0 1p

.Model Tranzistor NPN tr=5e-9 tf=8e-9

Vin in 0 pulse(0 5 0 1e-9 1e-9 1e-7 2e-7)
Vec ec 0 DC 5

[dc]
1
vin
0
5
0.1
[tran]
1e-9
6e-7
X
X
0
[ana]
1 2
0
1 1
1 1 0 5
3
v(in)
v(out)
v(ec)
0
1 1
1 1 0 5
2
v(in)
v(out)
[end]
