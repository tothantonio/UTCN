[aimspice]
[description]
264
Inversor NMOS static(analiza curent continuu)

!*Ordine parametri tranzistor NMOS: DGSB
M1 out in 0 0 NMOS1 l=1u w=1u
.Model NMOS1 nmos vto=1.5

M2 dd gg out out NMOS2 l=25u w=1u
.Model NMOS2 nmos vto=2.5

Vin in 0 DC 0
Vdd dd 0 DC 5
Vgg gg 0 DC 7.5


[dc]
1
Vin
0
5
0.1
[ana]
1 1
0
1 1
1 1 -1 6
2
v(out)
v(in)
[end]
