[aimspice]
[description]
390
Inversor NMOS static(analiza semnal pulse)

!*Ordinea parametrilor pentru tranzistorul NMOS: DGSB
M1 out in 0 0 NMOS1 l=1u w=1u
.Model NMOS1 nmos vto=1.5

M2 dd gg out out NMOS2 l=25u w=1u
.Model NMOS2 nmos vto=2.5

Vin in 0 pulse(0 5 0 1e-10 1e-10 1e-9 2e-9)
Vdd dd 0 DC 5
Vgg gg 0 DC 7.5

!*Vin=0V => M1 blocat => Vout=Vgg-Vt=7.5V-2.5V=5V
!*Vin=5V => M1 deschis => Vout=0V

[dc]
1
Vin
0
5
0.1
[tran]
1e-10
5e-9
X
X
0
[ana]
4 1
0
1 1
1 1 -1 6
2
v(out)
v(in)
[end]
