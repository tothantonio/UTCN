[aimspice]
[description]
326
Inversor cu tranzistor bipolar(analiza semnal pulse)
R1 in 1 1k
Rb 1 eb 7k
Rc out ec 1k
C1 in 1 30p

C2 0 out 1p
!*Acest condensator este pus ca sa corecteze iesirea inversorului

Q out 1 0 Tranzistor
.Model Tranzistor NPN tr=5e-9 tf=8e-9

Vin in 0 pulse(0 5 0 1e-9 1e-9 1e-7 2e-7)
Vec ec 0 DC 5
Veb eb 0 DC -1

[tran]
1e-9
5e-7
X
X
0
[ana]
4 1
0
1 1
1 1 -2 6
2
v(in)
v(out)
[end]
