[aimspice]
[description]
109
Redresor Monoalternanta
D1 1 2 diodaS
.Model diodaS D tt=1e-9
rl 2 0 100
vin 1 0 dc 5 sin(0 5 1k 0 0)


[tran]
1e-9
6e-3
0
0.0001
0
[ana]
4 1
0
1 1
1 1 -6 6
2
v(1)
v(2)
[end]
