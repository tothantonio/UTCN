[aimspice]
[description]
296
Stabilizator cu reac�ie f�r� amplificator de eroare
D1 1 2 dioda
D2 0 1 dioda
D3 0 3 dioda
D4 3 2 dioda
D5 0 Vz zener
C1 0 2 1m
R1 2 VZ 220
RL 0 out 100
Q1 2 Vz out tranzistor
Vin 1 3 sin(0 10 50 0 0)
.model dioda D TT=1e-9
.model zener D BV=6.8
.model tranzistor NPN tr=1e-9 tf=1e-9
[tran]
1e-9
60e-3
X
X
0
[ana]
4 1
0
1 1
1 1 -2 10
3
v(1)
v(outr)
v(2)
[end]
